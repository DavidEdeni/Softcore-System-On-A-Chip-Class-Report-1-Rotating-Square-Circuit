`timescale 1ns / 1ps // Defines this module's simulation time unit (1 ns) and time precision unit (1 ps)

module top( // Defines the top-level module for the overall circuit design of the Nexys4 DDR™ FPGA Board
    input logic CLK100MHZ, // Primary 100 MHz clock input signal from the FPGA board
    input logic [15:0] SW, // 16 input switch signals from the FPGA board
    output logic CA, // Output signal for the 'A' segment (cathode) of the 7-segment display
    output logic CB, // Output signal for the 'B' segment (cathode) of the 7-segment display
    output logic CC, // Output signal for the 'C' segment (cathode) of the 7-segment display
    output logic CD, // Output signal for the 'D' segment (cathode) of the 7-segment display
    output logic CE, // Output signal for the 'E' segment (cathode) of the 7-segment display
    output logic CF, // Output signal for the 'F' segment (cathode) of the 7-segment display
    output logic CG, // Output signal for the 'G' segment (cathode) of the 7-segment display
    output logic [7:0] An // 8 digit enable/Anode output signals for selecting which of the four-digit seven-segment display/8 7-segment digits is active
);

logic clk; // Internal, slower clock wire generated by the clockRate module
logic side; // Internal wire representing the "side" (half of rotation) for the digitSel module
logic [6:0] CX; // Internal wire for the 7-segment display pattern (segments A-G) for the segSel module

clockRate #(.N(29)) clockRate( // Instantiates the clockRate (counter) module with bit width parameter N = 29 (default value 29), this creates a 29-bit counter/clock
    .clk(CLK100MHZ), // Connect the 100 MHz input clock to the clockRate module
    .rst(0), // Connect a constant '0' for no reset (active high), rst = 0 → reset is off (the circuit runs normally)
    .en(1), // Connect a constant '1' to enable the clockRate (counter) module, en = 1 → clockRate (counter) is active
    .tic(clk) // Output the slower, divided clock tic to the internal "clk" wire
    );

digitSel digitSel( // Instantiates the digitSel module for 7-segment digit selection/multiplexing
    .En(SW[0]), // Connect input switch signal SW[0] as the Enable signal
    .Cw(SW[1]), // Connect input switch signal SW[1] as the Clockwise direction control
    .clk(clk), // Connect the slower, divided clock to the internal "clk" wire
    .side(side), // Output the "side" (top/bottom) signal to the internal "side" wire
    .An(An) // Output the 8-bit Anode selection to the Anode output signal pins
    );

segSel segSel( // Instantiates the segSel module for 7-segment pattern selection (segments A-G)
    .side(side), // Input the "side" (top/bottom) signal from the digitSel module
    .CX(CX) // Output the 7-bit segment pattern to the internal "CX" wire
    );
    
assign {CA, CB, CC, CD, CE, CF, CG} = CX[6:0]; // Assign the 7-bit segment pattern (CX) to the individual cathhode output pins (CA-CG)

endmodule // End of module definition